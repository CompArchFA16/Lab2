module fsm
(
	output misoBufe;
	output DMWriteEnable;
	output addressWriteEnable;
	output SRWriteEnable;
	output peripheralClkEdge;
	input shiftRegOutP;
	input conditioned;
);

endmodule